library verilog;
use verilog.vl_types.all;
entity MIPSGMN_vlg_vec_tst is
end MIPSGMN_vlg_vec_tst;
